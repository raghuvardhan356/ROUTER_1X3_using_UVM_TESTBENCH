package router_pkg;


//import uvm_pkg.sv
	import uvm_pkg::*;
//include uvm_macros.sv
	`include "uvm_macros.svh"
//`include "tb_defs.sv"
`include "src_xtn.sv"
`include "dst_xtn.sv"
`include "dst_sequence.sv"
`include "src_sequence.sv"
`include "src_agt_config.sv"
`include "dst_agt_config.sv"
`include "env_config.sv"
`include "src_sequencer.sv"
`include "src_driver.sv"
`include "src_monitor.sv"

`include "dst_sequencer.sv"
`include "dst_driver.sv"
`include "dst_monitor.sv"
`include "src_agt.sv"
`include "src_agt_top.sv"
//`include "ram_wr_seqs.sv"

//`include "read_xtn.sv"
//`include "dst_monitor.sv"
//`include "_driver.sv"
`include "dst_agt.sv"
`include "dst_agt_top.sv"

`include "virtual_sequencer.sv"
`include "virtual_sequence.sv"
`include "sb.sv"

`include "env.sv"


`include "router_test.sv"
endpackage
